// linear feedback shift registers to generate pseudorandom numbers
module lfsr(seed, value);
    input seed;
    
    output value;

endmodule
