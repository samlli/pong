module pong():



endmodule
