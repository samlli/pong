// outputs X and Y coordinates of upper left corner of paddle
module paddle(width, clk, reset, outX, outY, collision);



endmodule
